// stage_ex.v
// Execute stage
module stage_ex (
    input clk,
    input rst
);
    // ALU and execute logic
endmodule
