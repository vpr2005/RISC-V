// stage_wb.v
// Write-back stage
module stage_wb (
    input clk,
    input rst
);
    // Register file write-back
endmodule
