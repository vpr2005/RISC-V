// stage_mem.v
// Memory stage
module stage_mem (
    input clk,
    input rst
);
    // Data memory access
endmodule
