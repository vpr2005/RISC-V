// cpu_top.v
// Top-level module for 5-stage pipelined RISC-V processor

module cpu_top (
    input clk,
    input rst
);
    // Instantiate pipeline stages and hazard/forwarding units here
    // Connect pipeline registers and data paths
endmodule
